module hello_pli;
initial $hello;
endmodule
